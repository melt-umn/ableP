grammar edu:umn:cs:melt:ableP:extensions:syntax_check:ext ;

import edu:umn:cs:melt:ableP:concretesyntax ;

parser pp::Expr_c { edu:umn:cs:melt:ableP:extensions:tables ; }


