grammar edu:umn:cs:melt:ableP:host:extensions ;

exports edu:umn:cs:melt:ableP:host:extensions:embeddedC ;
exports edu:umn:cs:melt:ableP:host:extensions:v6 ;
exports edu:umn:cs:melt:ableP:host:extensions:typeChecking ;
