grammar edu:umn:cs:melt:ableP:host:core:abstractsyntax;

nonterminal Program with pp, errors, host<Program>, inlined<Program> ;

abstract production program
p::Program ::= u::Unit
{ production attribute newUnits::Unit with seqUnit ;
  newUnits := emptyUnit() ;
  forwards to programWithNewUnits( seqUnit(u, newUnits) ) ;
}

abstract production programWithNewUnits
p::Program ::= u::Unit
{ p.pp = "/* Promela code generated by ableP. */ \n\n" ++ u.pp ++
         "/* The end. */ \n" ;
  u.ppi = "" ;
  u.ppterm = "; \n" ;
  p.errors := u.errors;

  production attribute transformations :: [ Function(Program ::= Program) ]
    with ++ ;
  transformations := [ ] ; -- applyInRenameTransformation ] ;

  p.host = applyTransformations ( programWithNewUnits(u.host), transformations ) ;

--  p.host = applyInRenameTransformation (
--            programWithNewUnits(u.host) ) ;

  p.inlined = programWithNewUnits(u.inlined) ;

  u.env = emptyDefs();
  u.alluses = u.uses ;


  p.transformed = applyARewriteRule(p.rwrules_Program, p,
                    programWithNewUnits(u.transformed));
}

function applyTransformations
Program ::= p::Program trafos::[ Function(Program ::= Program) ] 
{ return
    if   null(trafos)
    then p
    else applyTransformations (  head(trafos)(p), tail(trafos) ) ;
}

