grammar edu:umn:cs:melt:ableP:terminals ;

terminal FOR_t 'for' lexer classes {promela,promela_kwd};
terminal IN_t 'in' ; -- lexer classes {promela,promela_kwd};
terminal DOTDOT_t '..' ;
