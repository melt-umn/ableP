grammar edu:umn:cs:melt:ableP:abstractsyntax ;

nonterminal Program ;
abstract production program 
p::Program ::= u::Units   { }

nonterminal Units ;
abstract production units_one
us::Units ::= u::Units { } 
abstract production units_snoc
us::Units ::= some::Units u::Unit { }

nonterminal Unit; 
