grammar edu:umn:cs:melt:ableP:host:core:coreParser ;

import edu:umn:cs:melt:ableP:host:core:concretesyntax
  only Program_c ;

parser promelaCoreParser :: Program_c {
 edu:umn:cs:melt:ableP:host:core:concretesyntax ;
}
