grammar edu:umn:cs:melt:ableP:extensions:syntax_check ;

import edu:umn:cs:melt:ableP:host:core:concretesyntax ;

parser extGrammar::Program_c { edu:umn:cs:melt:ableP:extensions:tables ; }

-- Maybe the type of extGrammar should be Expr_c ?

