grammar edu:umn:cs:melt:ableP:terminals ;

terminal FOR 'for' lexer classes {promela,promela_kwd};
terminal IN  'in' ; -- lexer classes {promela,promela_kwd};
terminal DOTDOT '..' ;
terminal SELECT 'select'   lexer classes {promela,promela_kwd};
