grammar edu:umn:cs:melt:ableP:host:extensions:v6 ;

terminal FOR 'for' lexer classes {promela,promela_kwd};
terminal IN  'in' ; -- lexer classes {promela,promela_kwd};
terminal DOTDOT '..' ;
terminal SELECT 'select'   lexer classes {promela,promela_kwd};
