grammar edu:umn:cs:melt:ableP:abstractsyntax;
import edu:umn:cs:melt:ableP:terminals;
