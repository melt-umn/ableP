grammar edu:umn:cs:melt:ableP:host:core ;

exports edu:umn:cs:melt:ableP:host:core:concretesyntax ;
exports edu:umn:cs:melt:ableP:host:core:abstractsyntax ;
exports edu:umn:cs:melt:ableP:host:core:terminals ;

exports edu:umn:cs:melt:ableP:host:core:coreParser ;

exports edu:umn:cs:melt:ableP:host:core:driver ;
