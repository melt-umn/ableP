grammar edu:umn:cs:melt:ableP:host ;

exports edu:umn:cs:melt:ableP:host:core:terminals ;
exports edu:umn:cs:melt:ableP:host:core:concretesyntax ;
exports edu:umn:cs:melt:ableP:host:core:abstractsyntax ;

exports edu:umn:cs:melt:ableP:host:hostParser ;

exports edu:umn:cs:melt:ableP:host:driver ;

-- extensions
exports edu:umn:cs:melt:ableP:host:extensions:embeddedC ;
exports edu:umn:cs:melt:ableP:host:extensions:typeChecking ;
exports edu:umn:cs:melt:ableP:host:extensions:v6 ;



-- Need to allow qualifications and renaming on exports.

exports edu:umn:cs:melt:ableC:concretesyntax ; -- as AbleC ;
