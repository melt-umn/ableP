grammar edu:umn:cs:melt:ableP:abstractsyntax;

