grammar edu:umn:cs:melt:ableP:host:hostParser ;

import edu:umn:cs:melt:ableP:concretesyntax
  only Program_c ;

parser promelaParser :: Program_c {
 edu:umn:cs:melt:ableP:terminals ;
 edu:umn:cs:melt:ableP:concretesyntax ;

 edu:umn:cs:melt:ableC:terminals ;
 edu:umn:cs:melt:ableC:concretesyntax ;
}
