grammar edu:umn:cs:melt:ableP:host:core:abstractsyntax;

import edu:umn:cs:melt:ableP:host:core:terminals;

nonterminal Program with pp, errors, host<Program>, inlined<Program> ;

abstract production program
p::Program ::= u::Unit
{ production attribute newUnits::Unit with seqUnit ;
  newUnits := emptyUnit() ;
  forwards to programWithNewUnits( seqUnit(u, newUnits) ) ;
}

abstract production programWithNewUnits
p::Program ::= u::Unit
{ p.pp = "/* Promela code generated by ableP. */ \n\n" ++ u.pp ++
         "/* The end. */ \n" ;
  u.ppi = "" ;
  u.ppterm = "; \n" ;
  p.errors := u.errors;
  p.host = programWithNewUnits(u.host);
  p.inlined = programWithNewUnits(u.inlined) ;

  u.env = emptyDefs();
  u.alluses = u.uses ;
}

