grammar edu:umn:cs:melt:ableP:host:core:concretesyntax ;
